`ifndef TOPLEVEL_PROBE_MONITOR_SV
`define TOPLEVEL_PROBE_MONITOR_SV

class toplevel_probe_monitor extends uvm_monitor;

  `uvm_component_utils(toplevel_probe_monitor)

  virtual toplevel_probe_if vif;

  toplevel_probe_config     m_config;

  uvm_analysis_port #(tx) analysis_port;

  tx m_trans;

  extern function new(string name, uvm_component parent);

  // Methods run_phase, and do_mon generated by setting monitor_inc in file ./toplevel_probe.tpl
  extern task run_phase(uvm_phase phase);
  // TODO
  // extern task do_mon();

endclass : toplevel_probe_monitor 


function toplevel_probe_monitor::new(string name, uvm_component parent);
  super.new(name, parent);
  analysis_port = new("analysis_port", this);
endfunction : new


task toplevel_probe_monitor::run_phase(uvm_phase phase);
  `uvm_info(get_type_name(), "run_phase", UVM_HIGH)

  m_trans = tx::type_id::create("m_trans");
  // do_mon();
endtask : run_phase


// Start of inlined include file generated_tb/tb/include/dummy.sv
// End of inlined include file

`endif // TOPLEVEL_PROBE_MONITOR_SV

