package verif_utils_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;

  `include "verif_utils_threads.sv"
  `include "verif_utils_delays.sv"

endpackage : verif_utils_pkg

