`ifndef FIFO_OUT_SEQUENCER_SV
`define FIFO_OUT_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(fifo_out_tx) fifo_out_sequencer_t;


`endif // FIFO_OUT_SEQUENCER_SV

