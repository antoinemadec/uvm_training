package top_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;

  import uvm_sw_ipc_pkg::*;

  `include "top_config.sv"
  `include "top_env.sv"

endpackage : top_pkg

