`ifndef UVM_SERVER_MONITOR_SV
`define UVM_SERVER_MONITOR_SV

class uvm_server_monitor extends uvm_monitor;

  `uvm_component_utils(uvm_server_monitor)

  virtual uvm_server_if vif;

  uvm_server_config     m_config;

  uvm_analysis_port #(uvm_server_tx) analysis_port;

  uvm_server_tx m_trans;
  uvm_server_tx m_trans_read;

  extern function new(string name, uvm_component parent);

  // Methods run_phase, and do_mon generated by setting monitor_inc in file ./uvm_server.tpl
  extern task run_phase(uvm_phase phase);
  extern task do_mon();

endclass : uvm_server_monitor 


function uvm_server_monitor::new(string name, uvm_component parent);
  super.new(name, parent);
  analysis_port = new("analysis_port", this);
endfunction : new


task uvm_server_monitor::run_phase(uvm_phase phase);
  `uvm_info(get_type_name(), "run_phase", UVM_HIGH)

  m_trans = uvm_server_tx::type_id::create("m_trans");
  m_trans_read = uvm_server_tx::type_id::create("m_trans_read");
  do_mon();
endtask : run_phase


task uvm_server_monitor::do_mon();
  wait(vif.cb.reset == 0);

  forever begin
    @(vif.cb);

    // prev cycle is a read cmd
    if (m_trans.rwb) begin
      m_trans_read.data = vif.cb.rdata;
      analysis_port.write(m_trans_read);
    end

    while (vif.cb.cen !== 1) begin
      @(vif.cb);
    end
    m_trans.addr = vif.cb.address;
    m_trans.rwb  = vif.cb.wen === 0;

    if (vif.cb.wen === 1) begin
      for (int i = 0; i < 4; i++) begin
        m_trans.data[i*8 +: 8] = vif.cb.wdata & {8{vif.cb.byteen[i]}};
      end
      analysis_port.write(m_trans);
    end
    else begin
      m_trans_read.copy(m_trans);
    end
  end
endtask : do_mon

`endif // UVM_SERVER_MONITOR_SV

