`ifndef TOPLEVEL_PROBE_SEQUENCER_SV
`define TOPLEVEL_PROBE_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(tx) toplevel_probe_sequencer_t;


`endif // TOPLEVEL_PROBE_SEQUENCER_SV

