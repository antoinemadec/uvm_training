package toplevel_probe_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;


  `include "toplevel_probe_tx.sv"
  `include "toplevel_probe_config.sv"
  `include "toplevel_probe_driver.sv"
  `include "toplevel_probe_monitor.sv"
  `include "toplevel_probe_sequencer.sv"
  `include "toplevel_probe_coverage.sv"
  `include "toplevel_probe_agent.sv"
  `include "toplevel_probe_seq_lib.sv"

endpackage : toplevel_probe_pkg
